`ifndef ${TOP_IF}_SV
`define ${TOP_IF}_SV

interface ${top_if}(input clk, input rstn);

    //IO HERE
    //logic ...

endinterface
`endif